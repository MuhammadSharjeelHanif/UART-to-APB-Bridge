interface the_inp_intf_apb (input clk);
	
	logic 			PREADY;
	logic [31:0] 	PRDATA;


endinterface : the_inp_intf_apb