interface the_out_intf_uart (input clk);
	
	logic 				tx;
	
endinterface : the_out_intf_uart