interface the_inp_intf_uart (input clk);
	
	logic 		rx;

endinterface : the_inp_intf_uart