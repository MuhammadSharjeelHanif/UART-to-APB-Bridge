class out_monitor_uart extends  uvm_monitor;
	`uvm_component_utils(out_monitor_uart)

	function new(string name = "out_monitor_uart", uvm_component parent=null);
		super.new(name, parent);
	endfunction : new

/*-------------------------------------------------------------------------------
-- Interface, port, fields
-------------------------------------------------------------------------------*/
  uvm_analysis_port#(seq_item_uart) mon_analysis_port;
  virtual the_out_intf_uart vif;
  int baud_delay = 868;
  
  seq_item_uart rec ;

/*-------------------------------------------------------------------------------
-- Functions
-------------------------------------------------------------------------------*/
  // =============================
  // Build Phase Method
  // =============================
	virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    if (!uvm_config_db#(virtual the_out_intf_uart)::get(this, "", "the_out_intf_uart", vif)) // getting  the value from tb
      `uvm_fatal("OUT_MONITOR_uart", "Could not get vif")

    mon_analysis_port = new ("mon_analysis_port", this);
  endfunction // build_phase


  // =============================
  // Main Phase Method
  // =============================
  virtual task main_phase(uvm_phase phase);
    super.main_phase(phase);
    fork
      collect_data();
    join_none
    
  endtask // main_phase

  // =============================
  // Collecting data
  // =============================
  task collect_data;
    bit [7:0] data;

  	forever begin
      @(posedge vif.clk);

  		if (!vif.tx) begin
        repeat(baud_delay + (baud_delay / 2)) @(posedge vif.clk);
        
        for (int i = 0; i < 8; i++) begin
          data[i] = vif.tx;
          repeat(baud_delay) @(posedge vif.clk);
        end

        rec = seq_item_uart::type_id::create("OUT Monitor Pkt");
  			rec.tx = data;
        mon_analysis_port.write(rec);
        rec.display_seq_item_uart("OUT_MONITOR_uart");  
  		end
  	end
  endtask
endclass : out_monitor_uart